module inv8(input [0:7]x, output [0:7]y);
assign y = ~x;
endmodule
